module	TOP(
	input	clk,
	input	DRY,
	input	ovr_in,
	input	signed	[13:0]	AD,
	output	ad_clk,
    output  tx,
);

wire	ovr_out;
assign	ad_clk = clk;





endmodule 
